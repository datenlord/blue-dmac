import PcieTypes::*;
import DmaTypes::*;

module mkDmaController#() (DmaController ifc);


endmodule